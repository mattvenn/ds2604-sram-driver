`define assert(signal, value) \
        if (signal !== value) begin \
            $display("ASSERTION FAILED in %m: signal != value"); \
            $finish; \
        end

`timescale 1ns/1ns
`default_nettype none
module test;

    reg [12:0] address = 0;
    reg [7:0] data_write = 0;
    wire [7:0] data_read;

    inout [7:0] data;

    assign data = !n_we ? data_write : 8'bz;

    reg n_ce1 = 0;
    reg n_we = 0;
    reg n_oe = 0;
    reg ce2 = 0;
 
    integer i;

    /* Make a reset that pulses once. */
    initial begin

        $dumpfile("test.vcd");
        $dumpvars(0,test);
        # 800
       
        // read first 255 addresses and check data is correct
        // data generated by gen_mem.py
        for( i = 13'd0; i <= 13'd255; i ++ ) begin
            address <= i;
            ce2 <= 1;
            n_ce1 <= 0;
            n_oe <= 0;
            n_we <= 1;
            # 250;
            `assert(data, i);
        end

        # 800

        // write first 255 addresses back to front
        for( i = 13'd0; i <= 13'd255; i ++ ) begin
            address <= i;
            data_write <= 8'd255 - i;
            ce2 <= 1;
            n_ce1 <= 0;
            n_oe <= 1;
            n_we <= 0;
            # 250;
        end

        # 800
        // read first 255 addresses and check data is correct
        // data written by routine above
        for( i = 13'd0; i <= 13'd255; i ++ ) begin
            address <= i;
            ce2 <= 1;
            n_ce1 <= 0;
            n_oe <= 0;
            n_we <= 1;
            # 250;
            `assert(data, 8'd255 - i);
        end

        $finish;

    end

    // about 12mhz with 1ns timescale
    reg clk = 0;
    always #80 clk = !clk;

    ds2064 ds2064_inst (.address(address), .data(data), .n_ce1(n_ce1), .ce2(ce2), .n_we(n_we), .n_oe(n_oe));

    endmodule
